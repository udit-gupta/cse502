module InstrnInfo(inst_info);
output logic[22:0] inst_info[255];

initial begin

// numop(2),op1(2),op2(2),sizeop1(2),sizeop2(2),op1regno(4),op2regnum(4), ...GRP(5)    
inst_info[0]   = 23'b10010000000000000000000; //ADD     " ;
inst_info[1]   = 23'b10010011110000000000000; //ADD     " ;
inst_info[2]   = 23'b10000100000000000000000; //ADD     " ;
inst_info[3]   = 23'b10000111110000000000000; //ADD     " ;
inst_info[4]   = 23'b10111000000000000000000; //ADD     " ;
inst_info[5]   = 23'b10111011100000000000000; //ADD     " ;
inst_info[6]   = 23'b00000000000000000000000; //PUSH    " ;
inst_info[7]   = 23'b00000000000000000000000; //POP     " ;
inst_info[8]   = 23'b10010000000000000000000; //OR      " ;
inst_info[9]   = 23'b10010011110000000000000; //OR      " ;
inst_info[10]  = 23'b10000100000000000000000; //OR      " ;
inst_info[11]  = 23'b10000111110000000000000; //OR      " ;
inst_info[12]  = 23'b10001000000000000000000; //OR      " ;
inst_info[13]  = 23'b10001011100000000000000; //OR      " ;
inst_info[14]  = 23'b00000000000000000000000; //PUSH    " ;
inst_info[15]  = 23'b10000111110000000000000; //ESC_OP  " ;
inst_info[16]  = 23'b00000000000000000000000; //ADC     " ;
inst_info[17]  = 23'b00000000000000000000000; //ADC     " ;
inst_info[18]  = 23'b00000000000000000000000; //ADC     " ;
inst_info[19]  = 23'b00000000000000000000000; //ADC     " ;
inst_info[20]  = 23'b00000000000000000000000; //ADC     " ;
inst_info[21]  = 23'b00000000000000000000000; //ADC     " ;
inst_info[22]  = 23'b00000000000000000000000; //PUSH    " ;
inst_info[23]  = 23'b00000000000000000000000; //POP     " ;
inst_info[24]  = 23'b00000000000000000000000; //SBB     " ;
inst_info[25]  = 23'b00000000000000000000000; //SBB     " ;
inst_info[26]  = 23'b00000000000000000000000; //SBB     " ;
inst_info[27]  = 23'b00000000000000000000000; //SBB     " ;
inst_info[28]  = 23'b00000000000000000000000; //SBB     " ;
inst_info[29]  = 23'b00000000000000000000000; //SBB     " ;
inst_info[30]  = 23'b00000000000000000000000; //PUSH    " ;
inst_info[31]  = 23'b00000000000000000000000; //POP     " ;
inst_info[32]  = 23'b10010000000000000000000; //AND     " ;
inst_info[33]  = 23'b10010011110000000000000; //AND     " ;
inst_info[34]  = 23'b10000100000000000000000; //AND     " ;
inst_info[35]  = 23'b10000111110000000000000; //AND     " ;
inst_info[36]  = 23'b10111000000000000000000; //AND     " ;  
inst_info[37]  = 23'b10111011100000000000000; //AND     " ;
inst_info[38]  = 23'b00000000000000000000000; //PFX_ES  " ;
inst_info[39]  = 23'b00000000000000000000000; //DAA     " ;
inst_info[40]  = 23'b00000000000000000000000; //SUB     " ;
inst_info[41]  = 23'b00000000000000000000000; //SUB     " ;
inst_info[42]  = 23'b00000000000000000000000; //SUB     " ;
inst_info[43]  = 23'b00000000000000000000000; //SUB     " ;
inst_info[44]  = 23'b00000000000000000000000; //SUB     " ;
inst_info[45]  = 23'b00000000000000000000000; //SUB     " ;
inst_info[46]  = 23'b00000000000000000000000; //PFX_CS  " ;
inst_info[47]  = 23'b00000000000000000000000; //DAS     " ;
inst_info[48]  = 23'b10010000000000000000000; //XOR     " ;
inst_info[49]  = 23'b10010011110000000000000; //XOR     " ;
inst_info[50]  = 23'b10000100000000000000000; //XOR     " ;
inst_info[51]  = 23'b10000111110000000000000; //XOR     " ;
inst_info[52]  = 23'b10111000000000000000000; //XOR     " ;
inst_info[53]  = 23'b10111011100000000000000; //XOR     " ;
inst_info[54]  = 23'b00000000000000000000000; //PFX_SS  " ;
inst_info[55]  = 23'b00000000000000000000000; //AAA     " ;
inst_info[56]  = 23'b00000000000000000000000; //CMP     " ;
inst_info[57]  = 23'b00000000000000000000000; //CMP     " ;
inst_info[58]  = 23'b00000000000000000000000; //CMP     " ;
inst_info[59]  = 23'b00000000000000000000000; //CMP     " ;
inst_info[60]  = 23'b00000000000000000000000; //CMP     " ;
inst_info[61]  = 23'b00000000000000000000000; //CMP     " ;
inst_info[62]  = 23'b00000000000000000000000; //PFX_DS  " ;
inst_info[63]  = 23'b00000000000000000000000; //AAS     " ;
inst_info[64]  = 23'b00000000000000000000000; //REX     " ;
inst_info[65]  = 23'b00000000000000000000000; //REX     " ;
inst_info[66]  = 23'b00000000000000000000000; //REX     " ;
inst_info[67]  = 23'b00000000000000000000000; //REX     " ;
inst_info[68]  = 23'b00000000000000000000000; //REX     " ;
inst_info[69]  = 23'b00000000000000000000000; //REX     " ;
inst_info[70]  = 23'b00000000000000000000000; //REX     " ;
inst_info[71]  = 23'b00000000000000000000000; //REX     " ;
inst_info[72]  = 23'b00000000000000000000000; //REX     " ;
inst_info[73]  = 23'b00000000000000000000000; //REX     " ;
inst_info[74]  = 23'b00000000000000000000000; //REX     " ;
inst_info[75]  = 23'b00000000000000000000000; //REX     " ;
inst_info[76]  = 23'b00000000000000000000000; //REX     " ;
inst_info[77]  = 23'b00000000000000000000000; //REX     " ;
inst_info[78]  = 23'b00000000000000000000000; //REX     " ;
inst_info[79]  = 23'b00000000000000000000000; //REX     " ;
inst_info[80]  = 23'b01110011000000000000000; //PUSH    " ;
inst_info[81]  = 23'b01110011000001000000000; //PUSH    " ;
inst_info[82]  = 23'b01110011000010000000000; //PUSH    " ;
inst_info[83]  = 23'b01110011000011000000000; //PUSH    " ;
inst_info[84]  = 23'b01110011000100000000000; //PUSH    " ;
inst_info[85]  = 23'b01110011000101000000000; //PUSH    " ;
inst_info[86]  = 23'b01110011000110000000000; //PUSH    " ;
inst_info[87]  = 23'b01110011000111000000000; //PUSH    " ;
inst_info[88]  = 23'b01110011000000000000000; //POP     " ;
inst_info[89]  = 23'b01110011000001000000000; //POP     " ;
inst_info[90]  = 23'b01110011000010000000000; //POP     " ;
inst_info[91]  = 23'b01110011000011000000000; //POP     " ;
inst_info[92]  = 23'b01110011000100000000000; //POP     " ;
inst_info[93]  = 23'b01110011000101000000000; //POP     " ;
inst_info[94]  = 23'b01110011000110000000000; //POP     " ;
inst_info[95]  = 23'b01110011000111000000000; //POP     " ;
inst_info[96]  = 23'b00000000000000000000000; //PUSHA   " ;
inst_info[97]  = 23'b00000000000000000000000; //POPA    " ;
inst_info[98]  = 23'b00000000000000000000000; //BOUND   " ;
inst_info[99]  = 23'b00000000000000000000000; //MOVSXD  " ;
inst_info[100] = 23'b00000000000000000000000; //PF_FS   " ;
inst_info[101] = 23'b00000000000000000000000; //PF_GS   " ;
inst_info[102] = 23'b00000000000000000000000; //PF_OP   " ;
inst_info[103] = 23'b00000000000000000000000; //PF_A    " ;
inst_info[104] = 23'b00000000000000000000000; //PUSH    " ;
inst_info[105] = 23'b00000000000000000000000; //IMUL    " ;
inst_info[106] = 23'b00000000000000000000000; //PUSH    " ;
inst_info[107] = 23'b00000000000000000000000; //IMUL    " ;
inst_info[108] = 23'b00000000000000000000000; //INS     " ;
inst_info[109] = 23'b00000000000000000000000; //INS     " ;
inst_info[110] = 23'b00000000000000000000000; //OUTS    " ;
inst_info[111] = 23'b00000000000000000000000; //OUTS    " ;
inst_info[112] = 23'b00000000000000000000000; //J       " ;
inst_info[113] = 23'b00000000000000000000000; //J       " ;
inst_info[114] = 23'b00000000000000000000000; //J       " ;
inst_info[115] = 23'b00000000000000000000000; //J       " ;
inst_info[116] = 23'b00000000000000000000000; //J       " ;
inst_info[117] = 23'b00000000000000000000000; //J       " ;
inst_info[118] = 23'b00000000000000000000000; //J       " ;
inst_info[119] = 23'b00000000000000000000000; //J       " ;
inst_info[120] = 23'b00000000000000000000000; //J       " ;
inst_info[121] = 23'b00000000000000000000000; //J       " ;
inst_info[122] = 23'b00000000000000000000000; //J       " ;
inst_info[123] = 23'b00000000000000000000000; //J       " ;
inst_info[124] = 23'b00000000000000000000000; //J       " ;
inst_info[125] = 23'b00000000000000000000000; //J       " ;
inst_info[126] = 23'b00000000000000000000000; //J       " ;
inst_info[127] = 23'b00000000000000000000000; //J       " ;
inst_info[128] = 23'b10011000000000000000000; //ADD/AND/XOR " ;
inst_info[129] = 23'b10011011100000000000000; //ADD/AND/XOR " ;
inst_info[130] = 23'b00000000000000000000000; //        " ;
inst_info[131] = 23'b10011011000000000000000; //ADD/AND/XOR " ;
inst_info[132] = 23'b00000000000000000000000; //TEST    " ;
inst_info[133] = 23'b00000000000000000000000; //TEST    " ;
inst_info[134] = 23'b00000000000000000000000; //XCHG    " ;
inst_info[135] = 23'b00000000000000000000000; //XCHG    " ;
inst_info[136] = 23'b10010000000000000000000; //MOV     " ;
inst_info[137] = 23'b10010011110000000000000; //MOV     " ;
inst_info[138] = 23'b10000100000000000000000; //MOV     " ;
inst_info[139] = 23'b10000111110000000000000; //MOV     " ;
inst_info[140] = 23'b10011100000000000000000; //MOV     " ;//*
inst_info[141] = 23'b00000000000000000000000; //LEA     " ;
inst_info[142] = 23'b10011100000000000000000; //MOV     " ;//*
inst_info[143] = 23'b00000000000000000000000; //POP     " ;
inst_info[144] = 23'b00000000000000000000000; //NOP     " ;
inst_info[145] = 23'b00000000000000000000000; //XCHG    " ;
inst_info[146] = 23'b00000000000000000000000; //XCHG    " ;
inst_info[147] = 23'b00000000000000000000000; //XCHG    " ;
inst_info[148] = 23'b00000000000000000000000; //XCHG    " ;
inst_info[149] = 23'b00000000000000000000000; //XCHG    " ;
inst_info[150] = 23'b00000000000000000000000; //XCHG    " ;
inst_info[151] = 23'b00000000000000000000000; //XCHG    " ;
inst_info[152] = 23'b00000000000000000000000; //CBW     " ;
inst_info[153] = 23'b00000000000000000000000; //CWD     " ;
inst_info[154] = 23'b00000000000000000000000; //CALL    " ;
inst_info[155] = 23'b00000000000000000000000; //WAIT    " ;
inst_info[156] = 23'b00000000000000000000000; //PUSHF   " ;
inst_info[157] = 23'b00000000000000000000000; //POPF    " ;
inst_info[158] = 23'b00000000000000000000000; //SAHF    " ;
inst_info[159] = 23'b00000000000000000000000; //LAHF    " ;
inst_info[160] = 23'b00000000000000000000000; //MOV     " ;//*
inst_info[161] = 23'b00000000000000000000000; //MOV     " ;//*
inst_info[162] = 23'b00000000000000000000000; //MOV     " ;//*
inst_info[163] = 23'b00000000000000000000000; //MOV     " ;//*
inst_info[164] = 23'b00000000000000000000000; //MOVS    " ;
inst_info[165] = 23'b00000000000000000000000; //MOVS    " ;
inst_info[166] = 23'b00000000000000000000000; //CMPS    " ;
inst_info[167] = 23'b00000000000000000000000; //CMPS    " ;
inst_info[168] = 23'b00000000000000000000000; //TEST    " ;
inst_info[169] = 23'b00000000000000000000000; //TEST    " ;
inst_info[170] = 23'b00000000000000000000000; //STOS    " ;
inst_info[171] = 23'b00000000000000000000000; //STOS    " ;
inst_info[172] = 23'b00000000000000000000000; //LODS    " ;
inst_info[173] = 23'b00000000000000000000000; //LODS    " ;
inst_info[174] = 23'b00000000000000000000000; //SCAS    " ;
inst_info[175] = 23'b00000000000000000000000; //SCAS    " ;
inst_info[176] = 23'b10001000000000000000000; //MOV    " ;
inst_info[177] = 23'b00000000000000000000000; //MOV     " ;
inst_info[178] = 23'b10000000000000000000000; //MOV     " ;
inst_info[179] = 23'b10000000000000000000000; //MOV     " ;
inst_info[180] = 23'b10000000000000000000000; //MOV     " ;
inst_info[181] = 23'b10000000000000000000000; //MOV     " ;
inst_info[182] = 23'b10000000000000000000000; //MOV     " ;
inst_info[183] = 23'b10000000000000000000000; //MOV     " ;
inst_info[184] = 23'b10001011110000000000000; //MOV     " ;
inst_info[185] = 23'b10111011110001000000000; //MOV     " ;
inst_info[186] = 23'b10111011110010000000000; //MOV     " ;
inst_info[187] = 23'b10111011110011000000000; //MOV     " ;
inst_info[188] = 23'b10111011110100000000000; //MOV     " ;
inst_info[189] = 23'b10111011110101000000000; //MOV     " ;
inst_info[190] = 23'b10111011110110000000000; //MOV     " ;
inst_info[191] = 23'b10111011110111000000000; //MOV     " ;
inst_info[192] = 23'b00000000000000000000000; //GRP2    " ;
inst_info[193] = 23'b00000000000000000000000; //GRP2    " ;
inst_info[194] = 23'b00000000000000000000000; //RET     " ;
inst_info[195] = 23'b00000000000000000000000; //RETQ    " ;
inst_info[196] = 23'b00000000000000000000000; //LES     " ;
inst_info[197] = 23'b00000000000000000000000; //LDS     " ;
inst_info[198] = 23'b10011000000000000000000; //MOV     " ;
inst_info[199] = 23'b10011011100000000000000; //MOV     " ;
inst_info[200] = 23'b00000000000000000000000; //ADD/AND " ;
inst_info[201] = 23'b00000000000000000000000; //ADD/AND " ;
inst_info[202] = 23'b00000000000000000000000; //RET     " ;
inst_info[203] = 23'b00000000000000000000000; //ADD/AND " ;
inst_info[204] = 23'b00000000000000000000000; //INT3    " ;
inst_info[205] = 23'b00000000000000000000000; //INT     " ;
inst_info[206] = 23'b00000000000000000000000; //INTO    " ;
inst_info[207] = 23'b00000000000000000000000; //IRET    " ;
inst_info[208] = 23'b00000000000000000000000; //SF_GRP2 " ;
inst_info[209] = 23'b00000000000000000000000; //SF_GRP2 " ;
inst_info[210] = 23'b00000000000000000000000; //SF_GRP2 " ;
inst_info[211] = 23'b00000000000000000000000; //SF_GRP2 " ;
inst_info[212] = 23'b00000000000000000000000; //AAM " ;
inst_info[213] = 23'b00000000000000000000000; // " ;
inst_info[214] = 23'b00000000000000000000000; //AAD " ;
inst_info[215] = 23'b00000000000000000000000; //XLAT    " ;
inst_info[216] = 23'b00000000000000000000000; //ESC     " ;
inst_info[217] = 23'b00000000000000000000000; //ESC     " ;
inst_info[218] = 23'b00000000000000000000000; //ESC     " ;
inst_info[219] = 23'b00000000000000000000000; //ESC     " ;
inst_info[220] = 23'b00000000000000000000000; //ESC     " ;
inst_info[221] = 23'b00000000000000000000000; //ESC     " ;
inst_info[222] = 23'b00000000000000000000000; //ESC     " ;
inst_info[223] = 23'b00000000000000000000000; //ESC     " ;
inst_info[224] = 23'b00000000000000000000000; //LOOPNE  " ;
inst_info[225] = 23'b00000000000000000000000; //LOOPE   " ;
inst_info[226] = 23'b00000000000000000000000; //LOOP    " ;
inst_info[227] = 23'b00000000000000000000000; //JRCXZ   " ;
inst_info[228] = 23'b00000000000000000000000; //IN      " ;
inst_info[229] = 23'b00000000000000000000000; //IN      " ;
inst_info[230] = 23'b00000000000000000000000; //OUT     " ;
inst_info[231] = 23'b00000000000000000000000; //OUT     " ;
inst_info[232] = 23'b01100010000000000000000; //CALL    " ;
inst_info[233] = 23'b00000000000000000000000; //JMP     " ;
inst_info[234] = 23'b00000000000000000000000; //JMP     " ;
inst_info[235] = 23'b01100000000000000000000; //JMP     " ;
inst_info[236] = 23'b00000000000000000000000; //IN      " ;
inst_info[237] = 23'b00000000000000000000000; //IN      " ;
inst_info[238] = 23'b00000000000000000000000; //OUT     " ;
inst_info[239] = 23'b00000000000000000000000; //OUT     " ;
inst_info[240] = 23'b00000000000000000000000; //LOCK    " ;//*
inst_info[241] = 23'b00000000000000000000000; //        " ;//*
inst_info[242] = 23'b00000000000000000000000; //REPNE   " ;//*
inst_info[243] = 23'b00000000000000000000000; //REPE    " ;//*
inst_info[244] = 23'b00000000000000000000000; //HLT     " ;*
inst_info[245] = 23'b00000000000000000000000; //CMC     " ;
inst_info[246] = 23'b01010000000000000000000; //IMUL    " ;
inst_info[247] = 23'b01010011000000000000000; //IMUL    " ;
inst_info[248] = 23'b00000000000000000000000; //CLC     " ;
inst_info[249] = 23'b00000000000000000000000; //STC     " ;
inst_info[250] = 23'b00000000000000000000000; //CLI     " ;
inst_info[251] = 23'b00000000000000000000000; //STI     " ;
inst_info[252] = 23'b00000000000000000000000; //CLD     " ;
inst_info[253] = 23'b00000000000000000000000; //STD     " ;
inst_info[254] = 23'b00000000000000000000000; //INC     " ;
inst_info[255] = 23'b00000000000000000000000; //DEC     " ;

if (inst_info[1] == 23'b 0 ); 

end
endmodule
