module InstrnInfo(inst_info);
output logic[23:0] inst_info[256];

initial begin

// assert(destreg==srcreg](1),numop(2),op1(2),op2(2),sizeop1(2),sizeop2(2),op1regno(4),op2regnum(4), ...GRP(5)    
inst_info[0]   = 24'b110010000000000000000000; //ADD     " ;
inst_info[1]   = 24'b110010011110000000000000; //ADD     " ;
inst_info[2]   = 24'b110000100000000000000000; //ADD     " ;
inst_info[3]   = 24'b110000111110000000000000; //ADD     " ;
inst_info[4]   = 24'b110111000000000000000000; //ADD     " ;
inst_info[5]   = 24'b110111011100000000000000; //ADD     " ;
inst_info[6]   = 24'b000000000000000000000000; //PUSH    " ;
inst_info[7]   = 24'b000000000000000000000000; //POP     " ;
inst_info[8]   = 24'b110010000000000000000000; //OR      " ;
inst_info[9]   = 24'b110010011110000000000000; //OR      " ;
inst_info[10]  = 24'b110000100000000000000000; //OR      " ;
inst_info[11]  = 24'b110000111110000000000000; //OR      " ;
inst_info[12]  = 24'b110001000000000000000000; //OR      " ;
inst_info[13]  = 24'b110111011100000000000000; //OR      " ;
inst_info[14]  = 24'b000000000000000000000000; //PUSH    " ;
inst_info[15]  = 24'b110000111110000000000000; //ESC_OP  " ;
inst_info[16]  = 24'b000000000000000000000000; //ADC     " ;
inst_info[17]  = 24'b000000000000000000000000; //ADC     " ;
inst_info[18]  = 24'b000000000000000000000000; //ADC     " ;
inst_info[19]  = 24'b000000000000000000000000; //ADC     " ;
inst_info[20]  = 24'b000000000000000000000000; //ADC     " ;
inst_info[21]  = 24'b000000000000000000000000; //ADC     " ;
inst_info[22]  = 24'b000000000000000000000000; //PUSH    " ;
inst_info[23]  = 24'b000000000000000000000000; //POP     " ;
inst_info[24]  = 24'b000000000000000000000000; //SBB     " ;
inst_info[25]  = 24'b000000000000000000000000; //SBB     " ;
inst_info[26]  = 24'b000000000000000000000000; //SBB     " ;
inst_info[27]  = 24'b000000000000000000000000; //SBB     " ;
inst_info[28]  = 24'b000000000000000000000000; //SBB     " ;
inst_info[29]  = 24'b000000000000000000000000; //SBB     " ;
inst_info[30]  = 24'b000000000000000000000000; //PUSH    " ;
inst_info[31]  = 24'b000000000000000000000000; //POP     " ;
inst_info[32]  = 24'b110010000000000000000000; //AND     " ;
inst_info[33]  = 24'b110010011110000000000000; //AND     " ;
inst_info[34]  = 24'b110000100000000000000000; //AND     " ;
inst_info[35]  = 24'b110000111110000000000000; //AND     " ;
inst_info[36]  = 24'b110111000000000000000000; //AND     " ;  
inst_info[37]  = 24'b110111011100000000000000; //AND     " ;
inst_info[38]  = 24'b000000000000000000000000; //PFX_ES  " ;
inst_info[39]  = 24'b000000000000000000000000; //DAA     " ;
inst_info[40]  = 24'b000000000000000000000000; //SUB     " ;
inst_info[41]  = 24'b000000000000000000000000; //SUB     " ;
inst_info[42]  = 24'b000000000000000000000000; //SUB     " ;
inst_info[43]  = 24'b000000000000000000000000; //SUB     " ;
inst_info[44]  = 24'b000000000000000000000000; //SUB     " ;
inst_info[45]  = 24'b000000000000000000000000; //SUB     " ;
inst_info[46]  = 24'b000000000000000000000000; //PFX_CS  " ;
inst_info[47]  = 24'b000000000000000000000000; //DAS     " ;
inst_info[48]  = 24'b110010000000000000000000; //XOR     " ;
inst_info[49]  = 24'b110010011110000000000000; //XOR     " ;
inst_info[50]  = 24'b110000100000000000000000; //XOR     " ;
inst_info[51]  = 24'b110000111110000000000000; //XOR     " ;
inst_info[52]  = 24'b110111000000000000000000; //XOR     " ;
inst_info[53]  = 24'b110111011100000000000000; //XOR     " ;
inst_info[54]  = 24'b000000000000000000000000; //PFX_SS  " ;
inst_info[55]  = 24'b000000000000000000000000; //AAA     " ;
inst_info[56]  = 24'b000000000000000000000000; //CMP     " ;
inst_info[57]  = 24'b000000000000000000000000; //CMP     " ;
inst_info[58]  = 24'b000000000000000000000000; //CMP     " ;
inst_info[59]  = 24'b000000000000000000000000; //CMP     " ;
inst_info[60]  = 24'b000000000000000000000000; //CMP     " ;
inst_info[61]  = 24'b000000000000000000000000; //CMP     " ;
inst_info[62]  = 24'b000000000000000000000000; //PFX_DS  " ;
inst_info[63]  = 24'b000000000000000000000000; //AAS     " ;
inst_info[64]  = 24'b000000000000000000000000; //REX     " ;
inst_info[65]  = 24'b000000000000000000000000; //REX     " ;
inst_info[66]  = 24'b000000000000000000000000; //REX     " ;
inst_info[67]  = 24'b000000000000000000000000; //REX     " ;
inst_info[68]  = 24'b000000000000000000000000; //REX     " ;
inst_info[69]  = 24'b000000000000000000000000; //REX     " ;
inst_info[70]  = 24'b000000000000000000000000; //REX     " ;
inst_info[71]  = 24'b000000000000000000000000; //REX     " ;
inst_info[72]  = 24'b000000000000000000000000; //REX     " ;
inst_info[73]  = 24'b000000000000000000000000; //REX     " ;
inst_info[74]  = 24'b000000000000000000000000; //REX     " ;
inst_info[75]  = 24'b000000000000000000000000; //REX     " ;
inst_info[76]  = 24'b000000000000000000000000; //REX     " ;
inst_info[77]  = 24'b000000000000000000000000; //REX     " ;
inst_info[78]  = 24'b000000000000000000000000; //REX     " ;
inst_info[79]  = 24'b000000000000000000000000; //REX     " ;
inst_info[80]  = 24'b001110011000000000000000; //PUSH    " ;
inst_info[81]  = 24'b001110011000001000000000; //PUSH    " ;
inst_info[82]  = 24'b001110011000010000000000; //PUSH    " ;
inst_info[83]  = 24'b001110011000011000000000; //PUSH    " ;
inst_info[84]  = 24'b001110011000100000000000; //PUSH    " ;
inst_info[85]  = 24'b001110011000101000000000; //PUSH    " ;
inst_info[86]  = 24'b001110011000110000000000; //PUSH    " ;
inst_info[87]  = 24'b001110011000111000000000; //PUSH    " ;
inst_info[88]  = 24'b001110011000000000000000; //POP     " ;
inst_info[89]  = 24'b001110011000001000000000; //POP     " ;
inst_info[90]  = 24'b001110011000010000000000; //POP     " ;
inst_info[91]  = 24'b001110011000011000000000; //POP     " ;
inst_info[92]  = 24'b001110011000100000000000; //POP     " ;
inst_info[93]  = 24'b001110011000101000000000; //POP     " ;
inst_info[94]  = 24'b001110011000110000000000; //POP     " ;
inst_info[95]  = 24'b001110011000111000000000; //POP     " ;
inst_info[96]  = 24'b000000000000000000000000; //PUSHA   " ;
inst_info[97]  = 24'b000000000000000000000000; //POPA    " ;
inst_info[98]  = 24'b000000000000000000000000; //BOUND   " ;
inst_info[99]  = 24'b000000000000000000000000; //MOVSXD  " ;
inst_info[100] = 24'b000000000000000000000000; //PF_FS   " ;
inst_info[101] = 24'b000000000000000000000000; //PF_GS   " ;
inst_info[102] = 24'b000000000000000000000000; //PF_OP   " ;
inst_info[103] = 24'b000000000000000000000000; //PF_A    " ;
inst_info[104] = 24'b000000000000000000000000; //PUSH    " ;
inst_info[105] = 24'b000000000000000000000000; //IMUL    " ;
inst_info[106] = 24'b000000000000000000000000; //PUSH    " ;
inst_info[107] = 24'b000000000000000000000000; //IMUL    " ;
inst_info[108] = 24'b000000000000000000000000; //INS     " ;
inst_info[109] = 24'b000000000000000000000000; //INS     " ;
inst_info[110] = 24'b000000000000000000000000; //OUTS    " ;
inst_info[111] = 24'b000000000000000000000000; //OUTS    " ;
inst_info[112] = 24'b000000000000000000000000; //J       " ;
inst_info[113] = 24'b000000000000000000000000; //J       " ;
inst_info[114] = 24'b000000000000000000000000; //J       " ;
inst_info[115] = 24'b000000000000000000000000; //J       " ;
inst_info[116] = 24'b000000000000000000000000; //J       " ;
inst_info[117] = 24'b000000000000000000000000; //J       " ;
inst_info[118] = 24'b000000000000000000000000; //J       " ;
inst_info[119] = 24'b000000000000000000000000; //J       " ;
inst_info[120] = 24'b000000000000000000000000; //J       " ;
inst_info[121] = 24'b000000000000000000000000; //J       " ;
inst_info[122] = 24'b000000000000000000000000; //J       " ;
inst_info[123] = 24'b000000000000000000000000; //J       " ;
inst_info[124] = 24'b000000000000000000000000; //J       " ;
inst_info[125] = 24'b000000000000000000000000; //J       " ;
inst_info[126] = 24'b000000000000000000000000; //J       " ;
inst_info[127] = 24'b000000000000000000000000; //J       " ;
inst_info[128] = 24'b110011000000000000000000; //ADD/AND/XOR " ;
inst_info[129] = 24'b110011011100000000000000; //ADD/AND/XOR " ;
inst_info[130] = 24'b000000000000000000000000; //        " ;
inst_info[131] = 24'b110011011000000000000000; //ADD/AND/XOR " ;
inst_info[132] = 24'b000000000000000000000000; //TEST    " ;
inst_info[133] = 24'b000000000000000000000000; //TEST    " ;
inst_info[134] = 24'b000000000000000000000000; //XCHG    " ;
inst_info[135] = 24'b000000000000000000000000; //XCHG    " ;
inst_info[136] = 24'b010010000000000000000000; //MOV     " ;
inst_info[137] = 24'b010010011110000000000000; //MOV     " ;
inst_info[138] = 24'b010000100000000000000000; //MOV     " ;
inst_info[139] = 24'b010000111110000000000000; //MOV     " ;
inst_info[140] = 24'b010011100000000000000000; //MOV     " ;//*
inst_info[141] = 24'b000000000000000000000000; //LEA     " ;
inst_info[142] = 24'b010011100000000000000000; //MOV     " ;//*
inst_info[143] = 24'b001010010000000000000000; //POP     " ;
inst_info[144] = 24'b000000000000000000000000; //NOP     " ;
inst_info[145] = 24'b000000000000000000000000; //XCHG    " ;
inst_info[146] = 24'b000000000000000000000000; //XCHG    " ;
inst_info[147] = 24'b000000000000000000000000; //XCHG    " ;
inst_info[148] = 24'b000000000000000000000000; //XCHG    " ;
inst_info[149] = 24'b000000000000000000000000; //XCHG    " ;
inst_info[150] = 24'b000000000000000000000000; //XCHG    " ;
inst_info[151] = 24'b000000000000000000000000; //XCHG    " ;
inst_info[152] = 24'b000000000000000000000000; //CBW     " ;
inst_info[153] = 24'b000000000000000000000000; //CWD     " ;
inst_info[154] = 24'b000000000000000000000000; //CALL    " ;
inst_info[155] = 24'b000000000000000000000000; //WAIT    " ;
inst_info[156] = 24'b000000000000000000000000; //PUSHF   " ;
inst_info[157] = 24'b000000000000000000000000; //POPF    " ;
inst_info[158] = 24'b000000000000000000000000; //SAHF    " ;
inst_info[159] = 24'b000000000000000000000000; //LAHF    " ;
inst_info[160] = 24'b000000000000000000000000; //MOV     " ;//*
inst_info[161] = 24'b000000000000000000000000; //MOV     " ;//*
inst_info[162] = 24'b000000000000000000000000; //MOV     " ;//*
inst_info[163] = 24'b000000000000000000000000; //MOV     " ;//*
inst_info[164] = 24'b000000000000000000000000; //MOVS    " ;
inst_info[165] = 24'b000000000000000000000000; //MOVS    " ;
inst_info[166] = 24'b000000000000000000000000; //CMPS    " ;
inst_info[167] = 24'b000000000000000000000000; //CMPS    " ;
inst_info[168] = 24'b000000000000000000000000; //TEST    " ;
inst_info[169] = 24'b000000000000000000000000; //TEST    " ;
inst_info[170] = 24'b000000000000000000000000; //STOS    " ;
inst_info[171] = 24'b000000000000000000000000; //STOS    " ;
inst_info[172] = 24'b000000000000000000000000; //LODS    " ;
inst_info[173] = 24'b000000000000000000000000; //LODS    " ;
inst_info[174] = 24'b000000000000000000000000; //SCAS    " ;
inst_info[175] = 24'b000000000000000000000000; //SCAS    " ;
inst_info[176] = 24'b010001000000000000000000; //MOV    " ;
inst_info[177] = 24'b000000000000000000000000; //MOV     " ;
inst_info[178] = 24'b010000000000000000000000; //MOV     " ;
inst_info[179] = 24'b010000000000000000000000; //MOV     " ;
inst_info[180] = 24'b010000000000000000000000; //MOV     " ;
inst_info[181] = 24'b010000000000000000000000; //MOV     " ;
inst_info[182] = 24'b010000000000000000000000; //MOV     " ;
inst_info[183] = 24'b010000000000000000000000; //MOV     " ;
inst_info[184] = 24'b010111011110000000000000; //MOV     " ;
inst_info[185] = 24'b010111011110001000000000; //MOV     " ;
inst_info[186] = 24'b010111011110010000000000; //MOV     " ;
inst_info[187] = 24'b010111011110011000000000; //MOV     " ;
inst_info[188] = 24'b010111011110100000000000; //MOV     " ;
inst_info[189] = 24'b010111011110101000000000; //MOV     " ;
inst_info[190] = 24'b010111011110110000000000; //MOV     " ;
inst_info[191] = 24'b010111011110111000000000; //MOV     " ;
inst_info[192] = 24'b000000000000000000000000; //GRP2    " ;
inst_info[193] = 24'b000000000000000000000000; //GRP2    " ;
inst_info[194] = 24'b000000000000000000000000; //RET     " ;
inst_info[195] = 24'b000000000000000000000000; //RETQ    " ;
inst_info[196] = 24'b000000000000000000000000; //LES     " ;
inst_info[197] = 24'b000000000000000000000000; //LDS     " ;
inst_info[198] = 24'b010011000000000000000000; //MOV     " ;
inst_info[199] = 24'b010011011100000000000000; //MOV     " ;
inst_info[200] = 24'b000000000000000000000000; //ADD/AND " ;
inst_info[201] = 24'b000000000000000000000000; //ADD/AND " ;
inst_info[202] = 24'b000000000000000000000000; //RET     " ;
inst_info[203] = 24'b000000000000000000000000; //ADD/AND " ;
inst_info[204] = 24'b000000000000000000000000; //INT3    " ;
inst_info[205] = 24'b000000000000000000000000; //INT     " ;
inst_info[206] = 24'b000000000000000000000000; //INTO    " ;
inst_info[207] = 24'b000000000000000000000000; //IRET    " ;
inst_info[208] = 24'b000000000000000000000000; //SF_GRP2 " ;
inst_info[209] = 24'b000000000000000000000000; //SF_GRP2 " ;
inst_info[210] = 24'b000000000000000000000000; //SF_GRP2 " ;
inst_info[211] = 24'b000000000000000000000000; //SF_GRP2 " ;
inst_info[212] = 24'b000000000000000000000000; //AAM " ;
inst_info[213] = 24'b000000000000000000000000; // " ;
inst_info[214] = 24'b000000000000000000000000; //AAD " ;
inst_info[215] = 24'b000000000000000000000000; //XLAT    " ;
inst_info[216] = 24'b000000000000000000000000; //ESC     " ;
inst_info[217] = 24'b000000000000000000000000; //ESC     " ;
inst_info[218] = 24'b000000000000000000000000; //ESC     " ;
inst_info[219] = 24'b000000000000000000000000; //ESC     " ;
inst_info[220] = 24'b000000000000000000000000; //ESC     " ;
inst_info[221] = 24'b000000000000000000000000; //ESC     " ;
inst_info[222] = 24'b000000000000000000000000; //ESC     " ;
inst_info[223] = 24'b000000000000000000000000; //ESC     " ;
inst_info[224] = 24'b000000000000000000000000; //LOOPNE  " ;
inst_info[225] = 24'b000000000000000000000000; //LOOPE   " ;
inst_info[226] = 24'b000000000000000000000000; //LOOP    " ;
inst_info[227] = 24'b000000000000000000000000; //JRCXZ   " ;
inst_info[228] = 24'b000000000000000000000000; //IN      " ;
inst_info[229] = 24'b000000000000000000000000; //IN      " ;
inst_info[230] = 24'b000000000000000000000000; //OUT     " ;
inst_info[231] = 24'b000000000000000000000000; //OUT     " ;
inst_info[232] = 24'b001100010000000000000000; //CALL    " ;
inst_info[233] = 24'b000000000000000000000000; //JMP     " ;
inst_info[234] = 24'b000000000000000000000000; //JMP     " ;
inst_info[235] = 24'b001100000000000000000000; //JMP     " ;
inst_info[236] = 24'b000000000000000000000000; //IN      " ;
inst_info[237] = 24'b000000000000000000000000; //IN      " ;
inst_info[238] = 24'b000000000000000000000000; //OUT     " ;
inst_info[239] = 24'b000000000000000000000000; //OUT     " ;
inst_info[240] = 24'b000000000000000000000000; //LOCK    " ;//*
inst_info[241] = 24'b000000000000000000000000; //        " ;//*
inst_info[242] = 24'b000000000000000000000000; //REPNE   " ;//*
inst_info[243] = 24'b000000000000000000000000; //REPE    " ;//*
inst_info[244] = 24'b000000000000000000000000; //HLT     " ;*
inst_info[245] = 24'b000000000000000000000000; //CMC     " ;
inst_info[246] = 24'b001010000000000000000000; //IMUL    " ;
inst_info[247] = 24'b001010011000000000000000; //IMUL    " ;
inst_info[248] = 24'b000000000000000000000000; //CLC     " ;
inst_info[249] = 24'b000000000000000000000000; //STC     " ;
inst_info[250] = 24'b000000000000000000000000; //CLI     " ;
inst_info[251] = 24'b000000000000000000000000; //STI     " ;
inst_info[252] = 24'b000000000000000000000000; //CLD     " ;
inst_info[253] = 24'b000000000000000000000000; //STD     " ;
inst_info[254] = 24'b000000000000000000000000; //INC     " ;
inst_info[255] = 24'b001010011000000000000000; //IMM_GRP!     " ;

if (inst_info[1] == 24'b0 ); 

end
endmodule
