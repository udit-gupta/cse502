module Opcodes2(op2,ModRM2);
typedef logic[63:0] mystring;
output mystring op2[0:255];
output logic[255:0] ModRM2 = 256'b0;

initial begin

	//opcode mnemonics;

op2[0] ="Grp6";
op2[1] ="Grp7";
op2[2] ="LAR";
op2[3] ="LSL";
op2[4] ="NULL";
op2[5] ="SYSCALL";
op2[6] ="CLTS";
op2[7] ="SYSRET";
op2[8] ="INVD";
op2[9] ="WBINVD";
op2[10] ="NULL";
op2[11] ="IOP2";
op2[12] ="NULL";
op2[13] ="pfw";
op2[14] ="NULL";
op2[15] ="NULL";
op2[16] ="VEC";
op2[17] ="VEC";
op2[18] ="VEC";
op2[19] ="VEC";
op2[20] ="VEC";
op2[21] ="VEC";
op2[22] ="VEC";
op2[23] ="VEC";
op2[24] ="pfgrp16";
op2[25] ="NULL";
op2[26] ="NULL";
op2[27] ="NULL";
op2[28] ="NULL";
op2[29] ="NULL";
op2[30] ="NULL";
op2[31] ="NOP";
op2[32] ="MOV";
op2[33] ="MOV";
op2[34] ="MOV";
op2[35] ="MOV";
op2[36] ="NULL";
op2[37] ="NULL";
op2[38] ="NULL";
op2[39] ="NULL";
op2[40] ="VEC";
op2[41] ="VEC";
op2[42] ="VEC";
op2[43] ="VEC";
op2[44] ="VEC";
op2[45] ="VEC";
op2[46] ="VEC";
op2[47] ="VEC";
op2[48] ="WRMSR";
op2[49] ="RDTSC";
op2[50] ="RDMSR";
op2[51] ="RDPMC";
op2[52] ="SYSENTER";
op2[53] ="SYSEXIT";
op2[54] ="NULL";
op2[55] ="GETSEC";
op2[56] ="ESC3";
op2[57] ="NULL";
op2[58] ="ESC3";
op2[59] ="NULL";
op2[60] ="NULL";
op2[61] ="NULL";
op2[62] ="NULL";
op2[63] ="NULL";
op2[64] ="CMOVcc";
op2[65] ="CMOVcc";
op2[66] ="CMOVcc";
op2[67] ="CMOVcc";
op2[68] ="CMOVcc";
op2[69] ="CMOVcc";
op2[70] ="CMOVcc";
op2[71] ="CMOVcc";
op2[72] ="CMOVcc";
op2[73] ="CMOVcc";
op2[74] ="CMOVcc";
op2[75] ="CMOVcc";
op2[76] ="CMOVcc";
op2[77] ="CMOVcc";
op2[78] ="CMOVcc";
op2[79] ="CMOVcc";
op2[80] ="VEC";
op2[81] ="VEC";
op2[82] ="VEC";
op2[83] ="VEC";
op2[84] ="VEC";
op2[85] ="VEC";
op2[86] ="VEC";
op2[87] ="VEC";
op2[88] ="VEC";
op2[89] ="VEC";
op2[90] ="VEC";
op2[91] ="VEC";
op2[92] ="VEC";
op2[93] ="VEC";
op2[94] ="VEC";
op2[95] ="VEC";
op2[96] ="VEC";
op2[97] ="VEC";
op2[98] ="VEC";
op2[99] ="VEC";
op2[100] ="VEC";
op2[101] ="VEC";
op2[102] ="VEC";
op2[103] ="VEC";
op2[104] ="VEC";
op2[105] ="VEC";
op2[106] ="VEC";
op2[107] ="VEC";
op2[108] ="VEC";
op2[109] ="VEC";
op2[110] ="movd";
op2[111] ="movq";
op2[112] ="VEC";
op2[113] ="VEC";
op2[114] ="VEC";
op2[115] ="VEC";
op2[116] ="VEC";
op2[117] ="VEC";
op2[118] ="VEC";
op2[119] ="VEC";
op2[120] ="VEC";
op2[121] ="VEC";
op2[122] ="VEC";
op2[123] ="VEC";
op2[124] ="VEC";
op2[125] ="VEC";
op2[126] ="movd";
op2[127] ="movq";
op2[128] ="J";
op2[129] ="J";
op2[130] ="J";
op2[131] ="J";
op2[132] ="J";
op2[133] ="J";
op2[134] ="J";
op2[135] ="J";
op2[136] ="J";
op2[137] ="J";
op2[138] ="J";
op2[139] ="J";
op2[140] ="J";
op2[141] ="J";
op2[142] ="J";
op2[143] ="J";
op2[144] ="SET";
op2[145] ="SET";
op2[146] ="SET";
op2[147] ="SET";
op2[148] ="SET";
op2[149] ="SET";
op2[150] ="SET";
op2[151] ="SET";
op2[152] ="SET";
op2[153] ="SET";
op2[154] ="SET";
op2[155] ="SET";
op2[156] ="SET";
op2[157] ="SET";
op2[158] ="SET";
op2[159] ="SET";
op2[160] ="PUSH";
op2[161] ="POP";
op2[162] ="CPUID";
op2[163] ="BT";
op2[164] ="SHLD";
op2[165] ="SHLD";
op2[166] ="NULL";
op2[167] ="NULL";
op2[168] ="PUSH";
op2[169] ="POP";
op2[170] ="RSM";
op2[171] ="BTS";
op2[172] ="SHRD";
op2[173] ="SHRD";
op2[174] ="Grp15";
op2[175] ="IMUL";
op2[176] ="CMPXCHG";
op2[177] ="CMPXCHG";
op2[178] ="LSS";
op2[179] ="BTR";
op2[180] ="LFS";
op2[181] ="LGS";
op2[182] ="MOVZX";
op2[183] ="MOVZX";
op2[184] ="JMPE";
op2[185] ="Grp10";
op2[186] ="Grp8";
op2[187] ="BTC";
op2[188] ="BSF";
op2[189] ="BSR";
op2[190] ="MOVSX";
op2[191] ="MOVSX";
op2[192] ="XADD";
op2[193] ="XADD";
op2[194] ="VEC";
op2[195] ="VEC";
op2[196] ="VEC";
op2[197] ="VEC";
op2[198] ="VEC";
op2[199] ="Grp9";
op2[200] ="BSWAP";
op2[201] ="BSWAP";
op2[202] ="BSWAP";
op2[203] ="BSWAP";
op2[204] ="BSWAP";
op2[205] ="BSWAP";
op2[206] ="BSWAP";
op2[207] ="BSWAP";
op2[208] ="VEC";
op2[209] ="VEC";
op2[210] ="VEC";
op2[211] ="VEC";
op2[212] ="VEC";
op2[213] ="VEC";
op2[214] ="VEC";
op2[215] ="VEC";
op2[216] ="VEC";
op2[217] ="VEC";
op2[218] ="VEC";
op2[219] ="VEC";
op2[220] ="VEC";
op2[221] ="VEC";
op2[222] ="VEC";
op2[223] ="VEC";
op2[224] ="VEC";
op2[225] ="VEC";
op2[226] ="VEC";
op2[227] ="VEC";
op2[228] ="VEC";
op2[229] ="VEC";
op2[230] ="VEC";
op2[231] ="VEC";
op2[232] ="VEC";
op2[233] ="VEC";
op2[234] ="VEC";
op2[235] ="VEC";
op2[236] ="VEC";
op2[237] ="VEC";
op2[238] ="VEC";
op2[239] ="VEC";
op2[240] ="VEC";
op2[241] ="VEC";
op2[242] ="VEC";
op2[243] ="VEC";
op2[244] ="VEC";
op2[245] ="VEC";
op2[246] ="VEC";
op2[247] ="VEC";
op2[248] ="VEC";
op2[249] ="VEC";
op2[250] ="VEC";
op2[251] ="VEC";
op2[252] ="VEC";
op2[253] ="VEC";
op2[254] ="VEC";
op2[255] ="NULL";

if (op2[1] == 0);
end

endmodule
